// 
// Designer: <student ID> 
//
module MAS_2input(
    input signed [4:0]Din1,
    input signed [4:0]Din2,
    input [1:0]Sel,
    input signed[4:0]Q,
    output [1:0]Tcmp,
    output signed reg [4:0]TDout,
    output signed reg [3:0]Dout
);

/*Write your design here*/

endmodule