// 
// Designer: P76111783
//
module Sbox(
    input [7:0] s,
    output reg [7:0] s_
    );

always @(s)
begin
    case (s)
        8'h00: s_=8'h63;
        8'h01: s_=8'h7c;
        8'h02: s_=8'h77;
        8'h03: s_=8'h7b;
        8'h04: s_=8'hf2;
        8'h05: s_=8'h6b;
        8'h06: s_=8'h6f;
        8'h07: s_=8'hc5;
        8'h08: s_=8'h30;
        8'h09: s_=8'h01;
        8'h0a: s_=8'h67;
        8'h0b: s_=8'h2b;
        8'h0c: s_=8'hfe;
        8'h0d: s_=8'hd7;
        8'h0e: s_=8'hab;
        8'h0f: s_=8'h76;
        8'h10: s_=8'hca;
        8'h11: s_=8'h82;
        8'h12: s_=8'hc9;
        8'h13: s_=8'h7d;
        8'h14: s_=8'hfa;
        8'h15: s_=8'h59;
        8'h16: s_=8'h47;
        8'h17: s_=8'hf0;
        8'h18: s_=8'had;
        8'h19: s_=8'hd4;
        8'h1a: s_=8'ha2;
        8'h1b: s_=8'haf;
        8'h1c: s_=8'h9c;
        8'h1d: s_=8'ha4;
        8'h1e: s_=8'h72;
        8'h1f: s_=8'hc0;
        8'h20: s_=8'hb7;
        8'h21: s_=8'hfd;
        8'h22: s_=8'h93;
        8'h23: s_=8'h26;
        8'h24: s_=8'h36;
        8'h25: s_=8'h3f;
        8'h26: s_=8'hf7;
        8'h27: s_=8'hcc;
        8'h28: s_=8'h34;
        8'h29: s_=8'ha5;
        8'h2a: s_=8'he5;
        8'h2b: s_=8'hf1;
        8'h2c: s_=8'h71;
        8'h2d: s_=8'hd8;
        8'h2e: s_=8'h31;
        8'h2f: s_=8'h15;
        8'h30: s_=8'h04;
        8'h31: s_=8'hc7;
        8'h32: s_=8'h23;
        8'h33: s_=8'hc3;
        8'h34: s_=8'h18;
        8'h35: s_=8'h96;
        8'h36: s_=8'h05;
        8'h37: s_=8'h9a;
        8'h38: s_=8'h07;
        8'h39: s_=8'h12;
        8'h3a: s_=8'h80;
        8'h3b: s_=8'he2;
        8'h3c: s_=8'heb;
        8'h3d: s_=8'h27;
        8'h3e: s_=8'hb2;
        8'h3f: s_=8'h75;
        8'h40: s_=8'h09;
        8'h41: s_=8'h83;
        8'h42: s_=8'h2c;
        8'h43: s_=8'h1a;
        8'h44: s_=8'h1b;
        8'h45: s_=8'h6e;
        8'h46: s_=8'h5a;
        8'h47: s_=8'ha0;
        8'h48: s_=8'h52;
        8'h49: s_=8'h3b;
        8'h4a: s_=8'hd6;
        8'h4b: s_=8'hb3;
        8'h4c: s_=8'h29;
        8'h4d: s_=8'he3;
        8'h4e: s_=8'h2f;
        8'h4f: s_=8'h84;
        8'h50: s_=8'h53;
        8'h51: s_=8'hd1;
        8'h52: s_=8'h00;
        8'h53: s_=8'hed;
        8'h54: s_=8'h20;
        8'h55: s_=8'hfc;
        8'h56: s_=8'hb1;
        8'h57: s_=8'h5b;
        8'h58: s_=8'h6a;
        8'h59: s_=8'hcb;
        8'h5a: s_=8'hbe;
        8'h5b: s_=8'h39;
        8'h5c: s_=8'h4a;
        8'h5d: s_=8'h4c;
        8'h5e: s_=8'h58;
        8'h5f: s_=8'hcf;
        8'h60: s_=8'hd0;
        8'h61: s_=8'hef;
        8'h62: s_=8'haa;
        8'h63: s_=8'hfb;
        8'h64: s_=8'h43;
        8'h65: s_=8'h4d;
        8'h66: s_=8'h33;
        8'h67: s_=8'h85;
        8'h68: s_=8'h45;
        8'h69: s_=8'hf9;
        8'h6a: s_=8'h02;
        8'h6b: s_=8'h7f;
        8'h6c: s_=8'h50;
        8'h6d: s_=8'h3c;
        8'h6e: s_=8'h9f;
        8'h6f: s_=8'ha8;
        8'h70: s_=8'h51;
        8'h71: s_=8'ha3;
        8'h72: s_=8'h40;
        8'h73: s_=8'h8f;
        8'h74: s_=8'h92;
        8'h75: s_=8'h9d;
        8'h76: s_=8'h38;
        8'h77: s_=8'hf5;
        8'h78: s_=8'hbc;
        8'h79: s_=8'hb6;
        8'h7a: s_=8'hda;
        8'h7b: s_=8'h21;
        8'h7c: s_=8'h10;
        8'h7d: s_=8'hff;
        8'h7e: s_=8'hf3;
        8'h7f: s_=8'hd2;
        8'h80: s_=8'hcd;
        8'h81: s_=8'h0c;
        8'h82: s_=8'h13;
        8'h83: s_=8'hec;
        8'h84: s_=8'h5f;
        8'h85: s_=8'h97;
        8'h86: s_=8'h44;
        8'h87: s_=8'h17;
        8'h88: s_=8'hc4;
        8'h89: s_=8'ha7;
        8'h8a: s_=8'h7e;
        8'h8b: s_=8'h3d;
        8'h8c: s_=8'h64;
        8'h8d: s_=8'h5d;
        8'h8e: s_=8'h19;
        8'h8f: s_=8'h73;
        8'h90: s_=8'h60;
        8'h91: s_=8'h81;
        8'h92: s_=8'h4f;
        8'h93: s_=8'hdc;
        8'h94: s_=8'h22;
        8'h95: s_=8'h2a;
        8'h96: s_=8'h90;
        8'h97: s_=8'h88;
        8'h98: s_=8'h46;
        8'h99: s_=8'hee;
        8'h9a: s_=8'hb8;
        8'h9b: s_=8'h14;
        8'h9c: s_=8'hde;
        8'h9d: s_=8'h5e;
        8'h9e: s_=8'h0b;
        8'h9f: s_=8'hdb;
        8'ha0: s_=8'he0;
        8'ha1: s_=8'h32;
        8'ha2: s_=8'h3a;
        8'ha3: s_=8'h0a;
        8'ha4: s_=8'h49;
        8'ha5: s_=8'h06;
        8'ha6: s_=8'h24;
        8'ha7: s_=8'h5c;
        8'ha8: s_=8'hc2;
        8'ha9: s_=8'hd3;
        8'haa: s_=8'hac;
        8'hab: s_=8'h62;
        8'hac: s_=8'h91;
        8'had: s_=8'h95;
        8'hae: s_=8'he4;
        8'haf: s_=8'h79;
        8'hb0: s_=8'he7;
        8'hb1: s_=8'hc8;
        8'hb2: s_=8'h37;
        8'hb3: s_=8'h6d;
        8'hb4: s_=8'h8d;
        8'hb5: s_=8'hd5;
        8'hb6: s_=8'h4e;
        8'hb7: s_=8'ha9;
        8'hb8: s_=8'h6c;
        8'hb9: s_=8'h56;
        8'hba: s_=8'hf4;
        8'hbb: s_=8'hea;
        8'hbc: s_=8'h65;
        8'hbd: s_=8'h7a;
        8'hbe: s_=8'hae;
        8'hbf: s_=8'h08;
        8'hc0: s_=8'hba;
        8'hc1: s_=8'h78;
        8'hc2: s_=8'h25;
        8'hc3: s_=8'h2e;
        8'hc4: s_=8'h1c;
        8'hc5: s_=8'ha6;
        8'hc6: s_=8'hb4;
        8'hc7: s_=8'hc6;
        8'hc8: s_=8'he8;
        8'hc9: s_=8'hdd;
        8'hca: s_=8'h74;
        8'hcb: s_=8'h1f;
        8'hcc: s_=8'h4b;
        8'hcd: s_=8'hbd;
        8'hce: s_=8'h8b;
        8'hcf: s_=8'h8a;
        8'hd0: s_=8'h70;
        8'hd1: s_=8'h3e;
        8'hd2: s_=8'hb5;
        8'hd3: s_=8'h66;
        8'hd4: s_=8'h48;
        8'hd5: s_=8'h03;
        8'hd6: s_=8'hf6;
        8'hd7: s_=8'h0e;
        8'hd8: s_=8'h61;
        8'hd9: s_=8'h35;
        8'hda: s_=8'h57;
        8'hdb: s_=8'hb9;
        8'hdc: s_=8'h86;
        8'hdd: s_=8'hc1;
        8'hde: s_=8'h1d;
        8'hdf: s_=8'h9e;
        8'he0: s_=8'he1;
        8'he1: s_=8'hf8;
        8'he2: s_=8'h98;
        8'he3: s_=8'h11;
        8'he4: s_=8'h69;
        8'he5: s_=8'hd9;
        8'he6: s_=8'h8e;
        8'he7: s_=8'h94;
        8'he8: s_=8'h9b;
        8'he9: s_=8'h1e;
        8'hea: s_=8'h87;
        8'heb: s_=8'he9;
        8'hec: s_=8'hce;
        8'hed: s_=8'h55;
        8'hee: s_=8'h28;
        8'hef: s_=8'hdf;
        8'hf0: s_=8'h8c;
        8'hf1: s_=8'ha1;
        8'hf2: s_=8'h89;
        8'hf3: s_=8'h0d;
        8'hf4: s_=8'hbf;
        8'hf5: s_=8'he6;
        8'hf6: s_=8'h42;
        8'hf7: s_=8'h68;
        8'hf8: s_=8'h41;
        8'hf9: s_=8'h99;
        8'hfa: s_=8'h2d;
        8'hfb: s_=8'h0f;
        8'hfc: s_=8'hb0;
        8'hfd: s_=8'h54;
        8'hfe: s_=8'hbb;
        8'hff: s_=8'h16;
    endcase
end
endmodule